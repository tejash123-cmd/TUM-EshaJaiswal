--------------------------------------------------------------------------------
-- Copyright 2021, Lehrstuhl für Rechnerarchitektur & Parallele Systeme,
-- Fakultät für Informatik, Technische Universität München
--------------------------------------------------------------------------------

--Libraries
library ieee;
use ieee.std_logic_1164.all;


entity rechner_tb is
end entity;

architecture test of rechner_tb is

    signal A,B : std_logic_vector(2 downto 0);
    signal SEL : std_logic;
    signal SEGMENTS_0, SEGMENTS_1 : std_logic_vector(6 downto 0);
begin
end architecture;
